module TwoBitShift(output data_out, input data_in);
	assign data_out = data_in << 2;
endmodule
