module ALUSelectTB()
	reg [3:0] FunctC,
	reg [31:0] A,B,
	wire [31:0] ALUOut,
	wire Zero);
	
	ALUSelect uut (.FucntC,.A,.B.ALUOut)
	
	initial begin 
	Assign A = 
	
	end
	
endmodule