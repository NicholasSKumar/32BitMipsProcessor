module ThirtyTwoBitMultiTB();
	reg [15:0] A;
	reg [15:0] B;
	wire [31:0] product;
	
	ThirtyTwoBitMulti uut(.A, .B,.product);
	initial begin
		
		A = 16'b1010101010101010;
		B = 16'b1010101010101010;
		//43690
		//43690
		//1908816100
		//01110001110001100011100011100100
		#20
		A = 16'b0010011100011010;
		B = 16'b0101110111000000;
		//10010
		//24000
		//240240000
		//1110010100011100010110000000
		#20
		A = 16'b0111010100110000;
		B = 16'b0110010001001000;
		//30000
		//24672
		//740160000
		//00101100000111011111001000000000
		#20
		B = 16'b0111010100110000;
		A = 16'b0110010001001000;
		//24672
		//30000
		//720160000
		//00101100000111011111001000000000
		#20
		A = 16'b1111111111111111;
		B = 16'b1111111111111111;
		//30000
		//24672
		//740160000
		//00101100000111011111001000000000
		
	
	end
endmodule 
