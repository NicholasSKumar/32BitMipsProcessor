module SixtyFourBitMulTB();
	reg [31:0] A;
	reg [31:0] B;
	wire [63:0] product;
	
	SixtyFourBitMul uut(.A, .B,.product);
	initial begin
		A = 17'b11010101010101010;
		B = 17'b01110010000111001;
		#5
		A = 32'b11100100001110011100111010000011;
		B = 32'b11000000111000110101101000110010;
		#5
		A = 32'b10010010100101110100110101100010;
		B = 32'b10001001001010100000101010000101;
		
		//43690
	
	end

endmodule